class rst_sqr extends uvm_sequencer #(rst_pkt);

  `uvm_component_utils(rst_sqr)

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

endclass