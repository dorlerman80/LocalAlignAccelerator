module SW_DUT #()
    (
        input logic clk,
        input logic rst_n
    );

endmodule